module inv_sqrt_lut (
    input  logic clk,
    input  logic [6:0]  addr,    
    output logic [15:0] slope,   
    output logic [15:0] base     
);
    always_ff @(posedge clk) begin
        case (addr)
            7'd0: begin slope <= 16'hFF01; base <= 16'hFFFF; end
            7'd1: begin slope <= 16'hFF04; base <= 16'hFF01; end
            7'd2: begin slope <= 16'hFF07; base <= 16'hFE06; end
            7'd3: begin slope <= 16'hFF0A; base <= 16'hFD0D; end
            7'd4: begin slope <= 16'hFF0D; base <= 16'hFC17; end
            7'd5: begin slope <= 16'hFF10; base <= 16'hFB24; end
            7'd6: begin slope <= 16'hFF12; base <= 16'hFA34; end
            7'd7: begin slope <= 16'hFF15; base <= 16'hF946; end
            7'd8: begin slope <= 16'hFF18; base <= 16'hF85B; end
            7'd9: begin slope <= 16'hFF1A; base <= 16'hF773; end
            7'd10: begin slope <= 16'hFF1D; base <= 16'hF68D; end
            7'd11: begin slope <= 16'hFF1F; base <= 16'hF5A9; end
            7'd12: begin slope <= 16'hFF21; base <= 16'hF4C8; end
            7'd13: begin slope <= 16'hFF24; base <= 16'hF3EA; end
            7'd14: begin slope <= 16'hFF26; base <= 16'hF30E; end
            7'd15: begin slope <= 16'hFF28; base <= 16'hF234; end
            7'd16: begin slope <= 16'hFF2B; base <= 16'hF15C; end
            7'd17: begin slope <= 16'hFF2D; base <= 16'hF087; end
            7'd18: begin slope <= 16'hFF2F; base <= 16'hEFB3; end
            7'd19: begin slope <= 16'hFF31; base <= 16'hEEE2; end
            7'd20: begin slope <= 16'hFF33; base <= 16'hEE13; end
            7'd21: begin slope <= 16'hFF35; base <= 16'hED46; end
            7'd22: begin slope <= 16'hFF37; base <= 16'hEC7C; end
            7'd23: begin slope <= 16'hFF39; base <= 16'hEBB3; end
            7'd24: begin slope <= 16'hFF3B; base <= 16'hEAEC; end
            7'd25: begin slope <= 16'hFF3D; base <= 16'hEA27; end
            7'd26: begin slope <= 16'hFF3F; base <= 16'hE964; end
            7'd27: begin slope <= 16'hFF41; base <= 16'hE8A3; end
            7'd28: begin slope <= 16'hFF43; base <= 16'hE7E4; end
            7'd29: begin slope <= 16'hFF44; base <= 16'hE727; end
            7'd30: begin slope <= 16'hFF46; base <= 16'hE66B; end
            7'd31: begin slope <= 16'hFF48; base <= 16'hE5B1; end
            7'd32: begin slope <= 16'hFF4A; base <= 16'hE4F9; end
            7'd33: begin slope <= 16'hFF4B; base <= 16'hE443; end
            7'd34: begin slope <= 16'hFF4D; base <= 16'hE38E; end
            7'd35: begin slope <= 16'hFF4F; base <= 16'hE2DB; end
            7'd36: begin slope <= 16'hFF50; base <= 16'hE22A; end
            7'd37: begin slope <= 16'hFF52; base <= 16'hE17A; end
            7'd38: begin slope <= 16'hFF53; base <= 16'hE0CC; end
            7'd39: begin slope <= 16'hFF55; base <= 16'hE020; end
            7'd40: begin slope <= 16'hFF57; base <= 16'hDF75; end
            7'd41: begin slope <= 16'hFF58; base <= 16'hDECB; end
            7'd42: begin slope <= 16'hFF59; base <= 16'hDE23; end
            7'd43: begin slope <= 16'hFF5B; base <= 16'hDD7C; end
            7'd44: begin slope <= 16'hFF5C; base <= 16'hDCD7; end
            7'd45: begin slope <= 16'hFF5E; base <= 16'hDC34; end
            7'd46: begin slope <= 16'hFF5F; base <= 16'hDB92; end
            7'd47: begin slope <= 16'hFF61; base <= 16'hDAF1; end
            7'd48: begin slope <= 16'hFF62; base <= 16'hDA51; end
            7'd49: begin slope <= 16'hFF63; base <= 16'hD9B3; end
            7'd50: begin slope <= 16'hFF65; base <= 16'hD916; end
            7'd51: begin slope <= 16'hFF66; base <= 16'hD87B; end
            7'd52: begin slope <= 16'hFF67; base <= 16'hD7E1; end
            7'd53: begin slope <= 16'hFF68; base <= 16'hD748; end
            7'd54: begin slope <= 16'hFF6A; base <= 16'hD6B0; end
            7'd55: begin slope <= 16'hFF6B; base <= 16'hD61A; end
            7'd56: begin slope <= 16'hFF6C; base <= 16'hD585; end
            7'd57: begin slope <= 16'hFF6D; base <= 16'hD4F1; end
            7'd58: begin slope <= 16'hFF6E; base <= 16'hD45E; end
            7'd59: begin slope <= 16'hFF70; base <= 16'hD3CD; end
            7'd60: begin slope <= 16'hFF71; base <= 16'hD33C; end
            7'd61: begin slope <= 16'hFF72; base <= 16'hD2AD; end
            7'd62: begin slope <= 16'hFF73; base <= 16'hD21F; end
            7'd63: begin slope <= 16'hFF74; base <= 16'hD192; end
            7'd64: begin slope <= 16'hFF75; base <= 16'hD106; end
            7'd65: begin slope <= 16'hFF76; base <= 16'hD07B; end
            7'd66: begin slope <= 16'hFF77; base <= 16'hCFF1; end
            7'd67: begin slope <= 16'hFF78; base <= 16'hCF69; end
            7'd68: begin slope <= 16'hFF79; base <= 16'hCEE1; end
            7'd69: begin slope <= 16'hFF7A; base <= 16'hCE5A; end
            7'd70: begin slope <= 16'hFF7B; base <= 16'hCDD5; end
            7'd71: begin slope <= 16'hFF7C; base <= 16'hCD50; end
            7'd72: begin slope <= 16'hFF7D; base <= 16'hCCCD; end
            7'd73: begin slope <= 16'hFF7E; base <= 16'hCC4A; end
            7'd74: begin slope <= 16'hFF7F; base <= 16'hCBC9; end
            7'd75: begin slope <= 16'hFF80; base <= 16'hCB48; end
            7'd76: begin slope <= 16'hFF81; base <= 16'hCAC8; end
            7'd77: begin slope <= 16'hFF82; base <= 16'hCA49; end
            7'd78: begin slope <= 16'hFF83; base <= 16'hC9CC; end
            7'd79: begin slope <= 16'hFF84; base <= 16'hC94F; end
            7'd80: begin slope <= 16'hFF85; base <= 16'hC8D3; end
            7'd81: begin slope <= 16'hFF86; base <= 16'hC858; end
            7'd82: begin slope <= 16'hFF87; base <= 16'hC7DD; end
            7'd83: begin slope <= 16'hFF87; base <= 16'hC764; end
            7'd84: begin slope <= 16'hFF88; base <= 16'hC6EB; end
            7'd85: begin slope <= 16'hFF89; base <= 16'hC674; end
            7'd86: begin slope <= 16'hFF8A; base <= 16'hC5FD; end
            7'd87: begin slope <= 16'hFF8B; base <= 16'hC587; end
            7'd88: begin slope <= 16'hFF8C; base <= 16'hC512; end
            7'd89: begin slope <= 16'hFF8C; base <= 16'hC49D; end
            7'd90: begin slope <= 16'hFF8D; base <= 16'hC42A; end
            7'd91: begin slope <= 16'hFF8E; base <= 16'hC3B7; end
            7'd92: begin slope <= 16'hFF8F; base <= 16'hC345; end
            7'd93: begin slope <= 16'hFF90; base <= 16'hC2D4; end
            7'd94: begin slope <= 16'hFF90; base <= 16'hC263; end
            7'd95: begin slope <= 16'hFF91; base <= 16'hC1F4; end
            7'd96: begin slope <= 16'hFF92; base <= 16'hC185; end
            7'd97: begin slope <= 16'hFF93; base <= 16'hC116; end
            7'd98: begin slope <= 16'hFF93; base <= 16'hC0A9; end
            7'd99: begin slope <= 16'hFF94; base <= 16'hC03C; end
            7'd100: begin slope <= 16'hFF95; base <= 16'hBFD0; end
            7'd101: begin slope <= 16'hFF95; base <= 16'hBF65; end
            7'd102: begin slope <= 16'hFF96; base <= 16'hBEFA; end
            7'd103: begin slope <= 16'hFF97; base <= 16'hBE90; end
            7'd104: begin slope <= 16'hFF97; base <= 16'hBE27; end
            7'd105: begin slope <= 16'hFF98; base <= 16'hBDBE; end
            7'd106: begin slope <= 16'hFF99; base <= 16'hBD56; end
            7'd107: begin slope <= 16'hFF99; base <= 16'hBCEF; end
            7'd108: begin slope <= 16'hFF9A; base <= 16'hBC89; end
            7'd109: begin slope <= 16'hFF9B; base <= 16'hBC23; end
            7'd110: begin slope <= 16'hFF9B; base <= 16'hBBBD; end
            7'd111: begin slope <= 16'hFF9C; base <= 16'hBB59; end
            7'd112: begin slope <= 16'hFF9D; base <= 16'hBAF5; end
            7'd113: begin slope <= 16'hFF9D; base <= 16'hBA91; end
            7'd114: begin slope <= 16'hFF9E; base <= 16'hBA2F; end
            7'd115: begin slope <= 16'hFF9E; base <= 16'hB9CC; end
            7'd116: begin slope <= 16'hFF9F; base <= 16'hB96B; end
            7'd117: begin slope <= 16'hFFA0; base <= 16'hB90A; end
            7'd118: begin slope <= 16'hFFA0; base <= 16'hB8A9; end
            7'd119: begin slope <= 16'hFFA1; base <= 16'hB84A; end
            7'd120: begin slope <= 16'hFFA1; base <= 16'hB7EA; end
            7'd121: begin slope <= 16'hFFA2; base <= 16'hB78C; end
            7'd122: begin slope <= 16'hFFA2; base <= 16'hB72E; end
            7'd123: begin slope <= 16'hFFA3; base <= 16'hB6D0; end
            7'd124: begin slope <= 16'hFFA4; base <= 16'hB673; end
            7'd125: begin slope <= 16'hFFA4; base <= 16'hB617; end
            7'd126: begin slope <= 16'hFFA5; base <= 16'hB5BB; end
            7'd127: begin slope <= 16'hFFA5; base <= 16'hB560; end
            default: begin slope <= 16'h0000; base <= 16'h0000; end
        endcase
    end

endmodule
